package async_fifo_pkg;

	`include "async_fifo_transaction.sv"
	`include "async_fifo_generator.sv"
	`include "async_fifo_driver.sv"
	`include "async_fifo_monitor.sv"
	`include "async_fifo_scoreboard.sv"
	`include "async_fifo_environment.sv"

endpackage
